`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:36:42 09/23/2019 
// Design Name: 
// Module Name:    comparador1b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module comparador1b(A,B,E,M);
xor(E,A,B)

if(A==1 && B==0)
M=1;
else
M=0;

endmodule
